`timescale 1ns / 1ps

//we're gonna have two clocks:
//a processing clock, at 50MHz (20ns)
//and a data clock, which is async
//(read from file) but which is at
//21.04MHz (47.53ns). how do you simulate that?
//
//so just getting data capture isn't going to be
//simulated here, since it's already done for you
//at this point in your saved data. we're going to
//have to address that at some point later on.
//(hint: you can cross clock domains with fifo_short_2clk)
//(generated by the fifo generator, but you can copy it)
//
//

//vsync module takes video from a monochrome camera
//with frame/line valid signals (like, say, a Quark)
//and outputs an AXI4 Stream Video compliant stream.
//this is synchronous to vclk so a downstream 2-clk
//FIFO handles that.
//
//ok let me think about this... the data is clocked in
//on the positive edge, which means we want to sample it
//on the negative edge. BUT we'd like all the subsequent
//blocks to use posedge, because AXI4-Stream is always
//sampled on the rising edge. we could just invert video_clk
//in the input buffer, before it gets wired anywhere.
//
//how do axi devices clock data out on the falling edge?
//i've never seen that. do we just depend on clock delay?
module vsync #(parameter WIDTH=8)
            (input vclk, //video clock
             input framevalid,
             input linevalid,
             input [WIDTH-1:0] data, //pixel data
             input reset, //AXI reset
             output [WIDTH-1:0] m_axis_data_tdata, //data output
             output m_axis_data_tlast,       //end of line
             input m_axis_data_tready,      //tready
             output m_axis_data_tvalid,      //tvalid
             output m_axis_data_tuser,       //start of frame
             output error);

   reg [WIDTH-1:0] data_flop;
   reg linevalid_flop, framevalid_flop, framevalid_flop_flop, sof_flop;

   wire vreset;

   reset_synchronizer inst_reset_synchronizer(
      .clk(vclk),
      .areset(reset),
      .reset(vreset)
   );

   wire eol;
   wire sof;

   always @(posedge vclk) begin
      if(vreset) begin
         data_flop <= 0;
         linevalid_flop <= 0;
         framevalid_flop <= 0;
         framevalid_flop_flop <= 0;
         sof_flop <= 0;
      end
      else begin
         data_flop <= data;
         linevalid_flop <= linevalid;
         framevalid_flop <= framevalid;
         framevalid_flop_flop <= framevalid_flop;
         sof_flop <= sof;
      end
   end

   assign eol = (~linevalid) & linevalid_flop;
   assign sof = linevalid & (~framevalid_flop_flop);

   assign m_axis_data_tdata = data_flop;
   assign m_axis_data_tlast = eol;
   assign m_axis_data_tvalid = (linevalid_flop & framevalid_flop);
   assign m_axis_data_tuser = sof_flop;
   assign error = 1'b0;

endmodule

