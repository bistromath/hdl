`timescale 1ns / 1ps

//we're gonna have two clocks:
//a processing clock, at 50MHz (20ns)
//and a data clock, which is async
//(read from file) but which is at
//21.04MHz (47.53ns). how do you simulate that?
//
//so just getting data capture isn't going to be
//simulated here, since it's already done for you
//at this point in your saved data. we're going to
//have to address that at some point later on.
//(hint: you can cross clock domains with fifo_short_2clk)
//(generated by the fifo generator, but you can copy it)
//
//

//vsync module takes video from a monochrome camera
//with frame/line valid signals (like, say, a Quark)
//and outputs an AXI4 Stream Video compliant stream.

module vsync #(parameter WIDTH=8)
            (input vclk, //video clock
             input framevalid,
             input linevalid,
             input [WIDTH-1:0] data, //pixel data
             input clk, //AXI clock
             input reset, //AXI reset
             output [WIDTH-1:0] m_axis_data_tdata, //data output
             output m_axis_data_tlast,       //end of line
             input m_axis_data_tready,      //tready
             output m_axis_data_tvalid,      //tvalid
             output m_axis_data_tuser,       //start of frame
             output error, //shit
             output overflow); //other shit

   reg [WIDTH-1:0] data_flop;
   reg linevalid_flop, framevalid_flop, framevalid_flop_flop, sof_flop;

   wire vreset;

   reset_synchronizer inst_reset_synchronizer(
      .clk(vclk),
      .areset(reset),
      .reset(vreset)
   );

   wire eol;
   wire sof;

   always @(posedge vclk) begin
      if(vreset) begin
         data_flop <= 0;
         linevalid_flop <= 0;
         framevalid_flop <= 0;
         framevalid_flop_flop <= 0;
         sof_flop <= 0;
      end
      else begin
         data_flop <= data;
         linevalid_flop <= linevalid;
         framevalid_flop <= framevalid;
         framevalid_flop_flop <= framevalid_flop;
         sof_flop <= sof;
      end
   end

   assign eol = (~linevalid) & linevalid_flop;
   assign sof = linevalid & (~framevalid_flop_flop);
   
   assign error = 0; //TODO: should do something with this.
   
   //1024-line 2-clock BRAM FIFO
   //input is non-flow-controlled,
   //so we just ignore the s_axis_tdata
   //and look for overflows.
   fifo_2clk_video inst_fifo_2clk_video(
      .s_aclk(vclk),
      .s_axis_tdata(data_flop),
      .s_axis_tlast(eol),
      .s_axis_tuser(sof_flop),
      .s_axis_tvalid(linevalid_flop & framevalid_flop),
      .s_axis_tready(), //we're always ready betch
      .m_aclk(clk),
      .s_aresetn(~reset),
      .m_axis_tdata(m_axis_data_tdata),
      .m_axis_tlast(m_axis_data_tlast),
      .m_axis_tuser(m_axis_data_tuser),
      .m_axis_tvalid(m_axis_data_tvalid),
      .m_axis_tready(m_axis_data_tready),
      .axis_overflow(overflow));
endmodule

